LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MultiPlexers IS
	GENERIC (
		REGISTER_SIZE : INTEGER
	);
	PORT (	
		D, R0, R1, R2, R3, R4, R5, R6, R7, G : IN STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		
		R_OUT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		D_OUT : IN STD_LOGIC;
		G_OUT : IN STD_LOGIC;
		
		BUS_OUT : OUT STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0)
	);
END MultiPlexers;

ARCHITECTURE dataflow OF MultiPlexers IS
BEGIN
	BUS_OUT <=
		D WHEN D_OUT='1' ELSE
		G WHEN G_OUT='1' ELSE
		R0 WHEN R_OUT(0) = '1' ELSE
		R1 WHEN R_OUT(1) = '1' ELSE
		R2 WHEN R_OUT(2) = '1' ELSE
		R3 WHEN R_OUT(3) = '1' ELSE
		R4 WHEN R_OUT(4) = '1' ELSE
		R5 WHEN R_OUT(5) = '1' ELSE
		R6 WHEN R_OUT(6) = '1' ELSE
		R7 WHEN R_OUT(7) = '1' ELSE
		(OTHERS => '0');
END dataflow;