LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ProgramCounter IS
	PORT (
		CLOCK : IN STD_LOGIC;
		CLEAR : IN STD_LOGIC;
		COUNT_NOW : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END ProgramCounter;

ARCHITECTURE behavior OF ProgramCounter IS
	SIGNAL COUNT : STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
	COUNT_NOW <= COUNT;

	PROCESS (CLOCK)
	BEGIN
		IF (RISING_EDGE(CLOCK)) THEN
			IF (CLEAR = '1') THEN
				COUNT <= "00";
			ELSE
				COUNT <= COUNT + 1;
			END IF;
		END IF;
	END PROCESS;
END behavior;
