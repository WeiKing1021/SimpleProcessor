LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY SimpleOp IS
	GENERIC (
		REGISTER_SIZE : INTEGER
	);
	PORT (
		OP_CODE : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		X_IN : IN STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		Y_IN : IN STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		OP_OUT : OUT STD_LOGIC_VECTOR(REGISTER_SIZE DOWNTO 0)
	);
END SimpleOp;

ARCHITECTURE dataflow OF SimpleOp IS
	SIGNAL X_NEW, Y_NEW : STD_LOGIC_VECTOR(REGISTER_SIZE DOWNTO 0);
BEGIN
	X_NEW <= '0' & X_IN;
	Y_NEW <= '0' & Y_IN;
	
	WITH OP_CODE SELECT OP_OUT <=
		X_NEW + Y_NEW WHEN "00",
		X_NEW - Y_NEW WHEN "01",
		X_NEW + 1 WHEN "10",
		X_NEW + 0 WHEN OTHERS;		
END dataflow;