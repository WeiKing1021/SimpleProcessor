-- LIBRARY
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- ENTITY AND PORT
ENTITY Dec4To16 IS
	PORT (
		ENABLE : IN STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END Dec4To16;

ARCHITECTURE dataflow OF Dec4To16 IS
BEGIN
	DATA_OUT <=
			"0000000000000000" WHEN ENABLE = '0' ELSE
			"0000000000000001" WHEN DATA_IN = "0000" ELSE
			"0000000000000010" WHEN DATA_IN = "0001" ELSE
			"0000000000000100" WHEN DATA_IN = "0010" ELSE
			"0000000000001000" WHEN DATA_IN = "0011" ELSE
			"0000000000010000" WHEN DATA_IN = "0100" ELSE
			"0000000000100000" WHEN DATA_IN = "0101" ELSE
			"0000000001000000" WHEN DATA_IN = "0110" ELSE
			"0000000010000000" WHEN DATA_IN = "0111" ELSE
			"0000000100000000" WHEN DATA_IN = "1000" ELSE
			"0000001000000000" WHEN DATA_IN = "1001" ELSE
			"0000010000000000" WHEN DATA_IN = "1010" ELSE
			"0000100000000000" WHEN DATA_IN = "1011" ELSE
			"0001000000000000" WHEN DATA_IN = "1100" ELSE
			"0010000000000000" WHEN DATA_IN = "1101" ELSE
			"0100000000000000" WHEN DATA_IN = "1110" ELSE
			"1000000000000000";			
END dataflow;