-- LIBRARY
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.all ;
USE IEEE.STD_LOGIC_SIGNED.ALL;

-- ENTITY AND PORT
ENTITY SimpleProcessor IS
	GENERIC (
		REGISTER_SIZE : INTEGER := 4
	);
	PORT (
		CLOCK : IN STD_LOGIC;
		ENABLE : IN STD_LOGIC;
		RESET : IN STD_LOGIC;

		DIN : IN STD_LOGIC_VECTOR(REGISTER_SIZE + 9 DOWNTO 0);

		REG0, REG1, REG2, REG3, REG4, REG5, REG6, REG7 : OUT STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		BUS_DATA : OUT STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		OVER_FLOW : OUT STD_LOGIC;
		DONE : OUT STD_LOGIC;
		STEP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END SimpleProcessor;

ARCHITECTURE behavior OF SimpleProcessor IS

	-- FLASH MEMORY
	COMPONENT MyRegister IS 
	GENERIC (
		REGISTER_SIZE : INTEGER
	);
	PORT (
		CLOCK : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		R_IN : IN STD_LOGIC; 
		DATA_OUT : OUT STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0)
	);
	END COMPONENT;
	
	-- DATA SELECTOR
	COMPONENT MultiPlexers IS
	GENERIC (
		REGISTER_SIZE : INTEGER
	);
	PORT (	
		D, R0, R1, R2, R3, R4, R5, R6, R7, G : IN STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		
		R_OUT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		D_OUT : IN STD_LOGIC;
		G_OUT : IN STD_LOGIC;
		
		BUS_OUT : OUT STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0)
	);
	END COMPONENT;
	
	-- ESSENTIAL PROCESS UNIT
	COMPONENT RealControlUnit IS
	GENERIC (
		REGISTER_SIZE : INTEGER
	);
	PORT (	
		CLOCK : IN STD_LOGIC;
		ENABLE : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		FUNCTION_IN : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		
		R_IN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		A_IN, G_IN : OUT STD_LOGIC;
		
		D_OUT : OUT STD_LOGIC;
		R_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		G_OUT : OUT STD_LOGIC;
		
		OP_CODE : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		
		PROCESS_DONE : OUT STD_LOGIC;
		PROCESS_STEP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);	
	END COMPONENT;
	
	-- SIMPLE OPERATOR
	COMPONENT SimpleOp IS
	GENERIC (
		REGISTER_SIZE : INTEGER
	);
	PORT (
		OP_CODE : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		X_IN : IN STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		Y_IN : IN STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
		OP_OUT : OUT STD_LOGIC_VECTOR(REGISTER_SIZE DOWNTO 0)
	);
	END COMPONENT;
		
	------------------
	-- SIGNAL START --
	------------------
	-- ESSENTIAL BUS SIGNAL
	SIGNAL DATA_BUS : STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
	
	
	-- FLUSH MEMORY IN GATE
	SIGNAL R_IN : STD_LOGIC_VECTOR(7 DOWNTO 0);
	
	-- A MEMORY IN GATE
	SIGNAL A_IN : STD_LOGIC;
	
	-- G MEMORY IN GATE
	SIGNAL G_IN : STD_LOGIC;
	
	
	-- FUNCTION DATA OUT GATE
	SIGNAL D_OUT : STD_LOGIC;
	
	-- FLUSH MEMORY OUT FATE
	SIGNAL R_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	
	-- G MEMORY OUT GATE
	SIGNAL G_OUT : STD_LOGIC;
	
	
	-- ALL BIT REGISTER
	SIGNAL D, R0, R1, R2, R3, R4, R5, R6, R7, G, A : STD_LOGIC_VECTOR(REGISTER_SIZE - 1 DOWNTO 0);
	
	
	-- OPERATOR TYPE CODE
	SIGNAL OP_CODE : STD_LOGIC_VECTOR(1 DOWNTO 0);
	
	-- OPERATOR RESULT SIGNAL
	SIGNAL OP_OUT : STD_LOGIC_VECTOR(REGISTER_SIZE DOWNTO 0);
BEGIN
	------------------
	-- REGISTER SET --
	------------------
	REG_0 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(0), R0);
	REG_1 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(1), R1);
	REG_2 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(2), R2);
	REG_3 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(3), R3);
	REG_4 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(4), R4);
	REG_5 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(5), R5);
	REG_6 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(6), R6);
	REG_7 : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, R_IN(7), R7);
	
	-- OTHER REGISTER
	REG_A : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (CLOCK, RESET, DATA_BUS, A_IN, A);
	REG_G : MyRegister GENERIC MAP (REGISTER_SIZE) PORT MAP (
		CLOCK, RESET, OP_OUT(REGISTER_SIZE - 1 DOWNTO 0), G_IN, G
	);
	
	-- MULTI PLEXER INSTANCE
	BUS_SELECTOR : MultiPlexers GENERIC MAP (REGISTER_SIZE) PORT MAP (
		D, R0, R1, R2, R3, R4, R5, R6, R7, G,
		R_OUT, D_OUT, G_OUT,
		DATA_BUS
	);
	
	-- OPERATOR INSTANCE
	OP : SimpleOp GENERIC MAP (REGISTER_SIZE) PORT MAP (OP_CODE, A, DATA_BUS, OP_OUT);
	
	-- ESSENTIAL CONTROL UNIT INSTANCE
	CONTROL_UNIT : RealControlUnit GENERIC MAP (REGISTER_SIZE) PORT MAP (
		CLOCK, ENABLE, RESET,
		DIN(REGISTER_SIZE + 9 DOWNTO REGISTER_SIZE + 0),
		R_IN, A_IN, G_IN,
		D_OUT, R_OUT, G_OUT,
		OP_CODE, DONE, STEP
	);
	
	-- D DATA
	D <= DIN(REGISTER_SIZE - 1 DOWNTO 0);
	
	-- OUTPUT
	REG0 <= R0;
	REG1 <= R1;
	REG2 <= R2;
	REG3 <= R3;
	REG4 <= R4;
	REG5 <= R5;
	REG6 <= R6;
	REG7 <= R7;
	
	-- BUS DATA
	BUS_DATA <= DATA_BUS;
	
	-- OPERATION OVERFLOW SIGNAL
	OVER_FLOW <= OP_OUT(REGISTER_SIZE);
END behavior;