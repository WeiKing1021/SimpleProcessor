LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY RealControlUnit IS
	GENERIC (
		REGISTER_SIZE : INTEGER
	);
	PORT (
		CLOCK : IN STD_LOGIC;
		ENABLE : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		FUNCTION_IN : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		
		R_IN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		A_IN, G_IN : OUT STD_LOGIC;
		
		D_OUT : OUT STD_LOGIC;
		R_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		G_OUT : OUT STD_LOGIC;
		
		OP_CODE : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		
		PROCESS_DONE : OUT STD_LOGIC;
		PROCESS_STEP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END RealControlUnit;

ARCHITECTURE dataflow OF RealControlUnit IS

	-- FUNCTION CACHE
	COMPONENT FunctionCache IS
	PORT (
		CLOCK : IN STD_LOGIC;
		FUNCTION_IN : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		FLUSH_FUNCTION : IN STD_LOGIC;
		FUNCTION_OUT : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
	END COMPONENT;
	
	-- PROGRAM COUNTER
	COMPONENT ProgramCounter IS
	PORT (
		CLOCK : IN STD_LOGIC;
		CLEAR : IN STD_LOGIC;
		COUNT_NOW : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
	END COMPONENT;
	
	-- 2 TO 4 DECODER
	COMPONENT Dec2To4 IS
	PORT (
		ENABLE : IN STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
	END COMPONENT;
	
	-- 3 TO 8 DECODER
	COMPONENT Dec3To8 IS
	PORT (
		ENABLE : IN STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
	END COMPONENT;
	
	-- 4 TO 16 DECODER
	COMPONENT Dec4To16 IS
	PORT (
		ENABLE : IN STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	END COMPONENT;
	
	------------------
	-- SIGNAL START --
	------------------
	
	-- FLUSH FUNCTION SIGNAL
	SIGNAL FLUSH_FUNCTION : STD_LOGIC;
	
	-- FUNCTION SIGNAL
	SIGNAL CACHE_FUNCTION, FINAL_FUNCTION : STD_LOGIC_VECTOR(9 DOWNTO 0);
	
	
	-- PROGRAM COUNTER CLEAR SIGNAL
	SIGNAL CLEAR : STD_LOGIC;
	-- PROGRAM COUNTER STEP
	SIGNAL STEP_NUM : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL STEP : STD_LOGIC_VECTOR(3 DOWNTO 0);
	-- PROCESS DOWN SIGNAL
	SIGNAL DONE : STD_LOGIC;
	
	
	-- FUNCTION SIGNAL
	SIGNAL COMMAND_NUM : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL X_NUM : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL Y_NUM : STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	-- DECODED FUNCTION SIGNAL
	SIGNAL COMMAND : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL X : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL Y : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	
	-- DETECT WHTHER CLEAR PROGRAM COUNTER
	CLEAR <= DONE OR (NOT(ENABLE) AND STEP(0));
	
	-- DETECT WHTHER ASSIGN NEW FUNCTION CACHE DATA
	FLUSH_FUNCTION <= ENABLE AND STEP(0);
	
	-- CHOOSE NEW FUNCTION OR CACHE FUNCTION
	FINAL_FUNCTION <= FUNCTION_IN WHEN STEP(0) = '1' ELSE CACHE_FUNCTION;
	
	-- SET COMMAND SIGNAL
	COMMAND_NUM <= FINAL_FUNCTION(9 DOWNTO 6);
	X_NUM <= FINAL_FUNCTION(5 DOWNTO 3);
	Y_NUM <= FINAL_FUNCTION(2 DOWNTO 0);
	
	-- DECODE COMMAND SIGNAL
	COMMAND_DECODER : Dec4To16 PORT MAP ('1', COMMAND_NUM, COMMAND);
	X_DECODER : Dec3To8 PORT MAP ('1', X_NUM, X);
	Y_DECODER : Dec3To8 PORT MAP ('1', Y_NUM, Y);
	
	-- FUNCTION CACHE INSTANCE
	FUNCTION_CACHE_ENTITY : FunctionCache
	PORT MAP (
		CLOCK,
		FUNCTION_IN,
		FLUSH_FUNCTION,
		CACHE_FUNCTION
	);
	
	-- PROGRAM COUNTER INSTANCE
	PRO_COUNTER : ProgramCounter PORT MAP (CLOCK, CLEAR, STEP_NUM);
	
	-- PROGRAM COUNTER DECODER
	COUNTER_DECODER : Dec2To4 PORT MAP ('1', STEP_NUM, STEP);
	
	-------------------
	-- BOOLEAN TABLE --
	-------------------
	R_IN_LOOP : FOR R IN 0 TO 7 GENERATE
		R_IN(R) <= 
			(COMMAND(0) AND STEP(0) AND X(R)) OR
			(COMMAND(1) AND STEP(0) AND X(R)) OR
			(COMMAND(2) AND STEP(2) AND X(R)) OR
			(COMMAND(3) AND STEP(2) AND X(R));
	END GENERATE R_IN_LOOP;
	
	R_OUT_LOOP : FOR R IN 0 TO 7 GENERATE
		R_OUT(R) <= 
			(COMMAND(0) AND STEP(0) AND Y(R)) OR
			-- COMMAND 2 NULL
			(COMMAND(2) AND STEP(0) AND X(R)) OR			
			(COMMAND(2) AND STEP(1) AND Y(R)) OR
			(COMMAND(3) AND STEP(0) AND X(R)) OR			
			(COMMAND(3) AND STEP(1) AND Y(R));
	END GENERATE R_OUT_LOOP;
	
	A_IN <= 
		(COMMAND(2) AND STEP(0)) OR
		(COMMAND(3) AND STEP(0));

	D_OUT <=
		(COMMAND(1) AND STEP(0));
		
	G_IN <=
		(COMMAND(2) AND STEP(1)) OR
		(COMMAND(3) AND STEP(1));
	
	G_OUT <=
		(COMMAND(2) AND STEP(2)) OR
		(COMMAND(3) AND STEP(2));
		
	OP_CODE <=
		"00" WHEN COMMAND(2) = '1' ELSE
		"01" WHEN COMMAND(3) = '1' ELSE
		"11";
		
	DONE <=
		(COMMAND(0) AND STEP(0)) OR
		(COMMAND(1) AND STEP(0)) OR
		(COMMAND(2) AND STEP(2)) OR
		(COMMAND(3) AND STEP(2));
		
	-- PROCESS STATE SYNC WITH CLOCK	
	PROCESS (CLOCK)
	BEGIN
		IF (RISING_EDGE(CLOCK)) THEN
			PROCESS_DONE <= DONE;
			PROCESS_STEP <= STEP_NUM;
		END IF;
	END PROCESS;
END dataflow;