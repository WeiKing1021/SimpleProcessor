LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY FunctionCache IS
	PORT (
		CLOCK : IN STD_LOGIC;
		FUNCTION_IN : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		FLUSH_FUNCTION : IN STD_LOGIC;
		FUNCTION_OUT : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END FunctionCache;

ARCHITECTURE behavior OF FunctionCache IS
	SIGNAL FUNCTION_CACHE : STD_LOGIC_VECTOR(9 DOWNTO 0);
BEGIN
	FUNCTION_OUT <= FUNCTION_CACHE;

	PROCESS (CLOCK)
	BEGIN
		IF (RISING_EDGE(CLOCK)) THEN
			IF (FLUSH_FUNCTION = '1') THEN
				FUNCTION_CACHE <= FUNCTION_IN;
			END IF;
		END IF;
	END PROCESS;
END behavior;